grammar edu:umn:cs:melt:exts:ableC:maps:src;

exports edu:umn:cs:melt:exts:ableC:maps:src:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:maps:src:concretesyntax;
