grammar edu:umn:cs:melt:exts:ableC:skeleton:src;

exports edu:umn:cs:melt:exts:ableC:skeleton:src:abstractsyntax;
exports edu:umn:cs:melt:exts:ableC:skeleton:src:concretesyntax;
