grammar edu:umn:cs:melt:exts:ableC:maps:src;

exports edu:umn:cs:melt:exts:ableC:maps:src:concretesyntax:typeExpr;
exports edu:umn:cs:melt:exts:ableC:maps:src:concretesyntax:constructor;
exports edu:umn:cs:melt:exts:ableC:maps:src:abstractsyntax;
